library verilog;
use verilog.vl_types.all;
entity tb_sha256 is
    generic(
        DEBUG           : integer := 0;
        CLK_HALF_PERIOD : integer := 2;
        CLK_PERIOD      : vl_notype;
        ADDR_NAME0      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_NAME1      : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        ADDR_VERSION    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        ADDR_CTRL       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        CTRL_INIT_VALUE : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        CTRL_NEXT_VALUE : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        CTRL_MODE_VALUE : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        ADDR_STATUS     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        STATUS_READY_BIT: integer := 0;
        STATUS_VALID_BIT: integer := 1;
        ADDR_BLOCK0     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        ADDR_BLOCK1     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        ADDR_BLOCK2     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        ADDR_BLOCK3     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        ADDR_BLOCK4     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        ADDR_BLOCK5     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        ADDR_BLOCK6     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        ADDR_BLOCK7     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        ADDR_BLOCK8     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        ADDR_BLOCK9     : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        ADDR_BLOCK10    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        ADDR_BLOCK11    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        ADDR_BLOCK12    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        ADDR_BLOCK13    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        ADDR_BLOCK14    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        ADDR_BLOCK15    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        ADDR_DIGEST0    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR_DIGEST1    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        ADDR_DIGEST2    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        ADDR_DIGEST3    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        ADDR_DIGEST4    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        ADDR_DIGEST5    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        ADDR_DIGEST6    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        ADDR_DIGEST7    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        SHA256_MODE     : integer := 1
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DEBUG : constant is 1;
    attribute mti_svvh_generic_type of CLK_HALF_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of CLK_PERIOD : constant is 3;
    attribute mti_svvh_generic_type of ADDR_NAME0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_NAME1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_VERSION : constant is 1;
    attribute mti_svvh_generic_type of ADDR_CTRL : constant is 1;
    attribute mti_svvh_generic_type of CTRL_INIT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of CTRL_NEXT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of CTRL_MODE_VALUE : constant is 1;
    attribute mti_svvh_generic_type of ADDR_STATUS : constant is 1;
    attribute mti_svvh_generic_type of STATUS_READY_BIT : constant is 1;
    attribute mti_svvh_generic_type of STATUS_VALID_BIT : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK2 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK3 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK4 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK5 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK6 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK7 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK8 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK9 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK10 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK11 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK12 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK13 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK14 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BLOCK15 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST0 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST1 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST2 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST3 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST4 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST5 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST6 : constant is 1;
    attribute mti_svvh_generic_type of ADDR_DIGEST7 : constant is 1;
    attribute mti_svvh_generic_type of SHA256_MODE : constant is 1;
end tb_sha256;
